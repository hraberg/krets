NON-LINEAR_DC_CKT.CIR - SIMPLE NON-LINEAR CIRCUIT
*
IS	0	1	DC	0.1A
*
R1	1	0	100
R2	1	2	10K
D1	2	0	DNOM
*
.MODEL DNOM D(IS=1E-15)
*
* ANALYSIS
.TRAN 	1MS  10MS
* VIEW RESULTS
.PRINT	TRAN 	V(1) V(2)
.PROBE
.END