Inverting opamp
v1 2 0 dc
e 3 0 0 one 999k
r1 3 one 3.29k
r2 one 2 1.18k
.dc v1 0 3.5 0.05
.print dc v(3,0)
.end