LINEAR_DC_CKT.CIR - SIMPLE CIRCUIT FOR NODAL ANALYSIS
*
IS	0	1	DC	1A
*
R1	1	0	10
R2	1	2	1K
R3	2	0	1K
*
* ANALYSIS
.TRAN 	1MS  10MS
* VIEW RESULTS
.PRINT	TRAN 	V(1) V(2)
.PROBE
.END