TRANSIENT_DC_CKT.CIR - SIMPLE CIRCUIT FOR TRANSIENT NODAL ANALYSIS
*
IS      0       1       DC      10A
*
R1      0       1       1
R2      1       2       1K
R3      2       0       100K
*
C1      0       2       10u
*
* ANALYSIS
.TRAN   0.0005 0.200
* VIEW RESULTS
.PLOT  TRAN    V(1) V(2)
* .PRINT  TRAN    V(1) V(2)
.PROBE
.END